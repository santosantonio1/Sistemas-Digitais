-- Registrador em que A=input, B=A, C=B, ...